library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prom_ic23 is
port (
	clk  : in  std_logic;
	ce   : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prom_ic23 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"04",X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"20",X"00",X"0C",X"0C",X"00",X"00",X"00",X"20",X"70",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"08",X"08",X"3E",X"08",X"08",X"00",X"10",X"10",X"10",X"FE",X"10",X"10",X"10",X"00",
		X"00",X"44",X"00",X"00",X"20",X"00",X"02",X"00",X"10",X"00",X"40",X"08",X"02",X"80",X"04",X"00",
		X"01",X"40",X"04",X"10",X"82",X"04",X"50",X"02",X"82",X"48",X"02",X"A0",X"08",X"45",X"20",X"02",
		X"3C",X"7E",X"DF",X"AF",X"D7",X"AF",X"56",X"3C",X"3C",X"42",X"99",X"BD",X"BD",X"99",X"42",X"3C",
		X"88",X"20",X"04",X"90",X"2A",X"56",X"0F",X"03",X"24",X"18",X"65",X"9A",X"1D",X"A0",X"56",X"28",
		X"3C",X"5A",X"AB",X"AD",X"D5",X"D3",X"6A",X"3C",X"38",X"68",X"DC",X"FA",X"2E",X"3F",X"16",X"0C",
		X"01",X"2A",X"54",X"2A",X"54",X"2A",X"54",X"80",X"3C",X"46",X"F9",X"8F",X"F3",X"9D",X"62",X"3C",
		X"08",X"08",X"1C",X"7F",X"1C",X"08",X"08",X"00",X"1C",X"3A",X"6D",X"75",X"77",X"36",X"1C",X"00",
		X"00",X"18",X"3C",X"7E",X"7E",X"3C",X"18",X"00",X"38",X"50",X"E8",X"F8",X"F0",X"D8",X"60",X"38",
		X"08",X"2A",X"1C",X"7F",X"1C",X"2A",X"08",X"00",X"38",X"4C",X"9D",X"BD",X"BD",X"B9",X"32",X"1C",
		X"62",X"91",X"09",X"3A",X"5C",X"90",X"89",X"46",X"3C",X"5E",X"EB",X"FF",X"DF",X"F7",X"7E",X"3C",
		X"FE",X"FC",X"F8",X"C0",X"80",X"10",X"60",X"80",X"F0",X"1C",X"06",X"83",X"C3",X"E3",X"F7",X"FE",
		X"FF",X"FF",X"BB",X"EE",X"EE",X"BC",X"F8",X"E0",X"E0",X"F8",X"FC",X"F6",X"BE",X"FF",X"6F",X"6B",
		X"40",X"10",X"80",X"C0",X"00",X"00",X"00",X"00",X"21",X"88",X"22",X"10",X"84",X"21",X"88",X"54",
		X"E5",X"D0",X"85",X"20",X"94",X"40",X"01",X"A0",X"40",X"10",X"44",X"90",X"02",X"A8",X"C5",X"E8",
		X"C0",X"E8",X"60",X"14",X"48",X"04",X"2A",X"01",X"00",X"00",X"80",X"28",X"40",X"10",X"C0",X"D0",
		X"FC",X"FC",X"F8",X"FC",X"F2",X"D9",X"0F",X"07",X"00",X"00",X"C0",X"C0",X"98",X"38",X"7C",X"FC",
		X"BB",X"D6",X"77",X"E6",X"8E",X"3C",X"F8",X"E0",X"E0",X"F8",X"3C",X"8E",X"66",X"F7",X"F6",X"EB",
		X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"03",X"05",X"0A",X"D4",X"E8",X"D0",X"B8",X"78",
		X"7F",X"EF",X"C7",X"C3",X"41",X"60",X"30",X"0F",X"01",X"06",X"08",X"01",X"03",X"1F",X"3F",X"7F",
		X"E7",X"E4",X"FC",X"7F",X"77",X"37",X"1E",X"07",X"07",X"1F",X"3D",X"7E",X"5E",X"FB",X"BE",X"BE",
		X"19",X"16",X"28",X"76",X"7B",X"FC",X"F8",X"E0",X"00",X"00",X"00",X"00",X"02",X"02",X"0C",X"0A",
		X"27",X"93",X"29",X"44",X"12",X"24",X"09",X"02",X"05",X"10",X"01",X"44",X"12",X"89",X"23",X"97",
		X"03",X"0B",X"10",X"05",X"12",X"00",X"00",X"00",X"80",X"48",X"20",X"15",X"28",X"06",X"27",X"13",
		X"39",X"33",X"07",X"0F",X"0F",X"03",X"00",X"00",X"E0",X"D0",X"CB",X"6F",X"3F",X"1F",X"3E",X"3C",
		X"DF",X"CB",X"ED",X"67",X"71",X"3C",X"1F",X"07",X"07",X"1F",X"3C",X"71",X"67",X"ED",X"CF",X"DA",
		X"1E",X"1D",X"0B",X"17",X"2B",X"50",X"A0",X"C0",X"00",X"00",X"00",X"03",X"07",X"0F",X"1F",X"1F",
		X"20",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"77",X"22",X"77",X"22",X"77",
		X"77",X"22",X"77",X"22",X"F7",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"20",
		X"F0",X"07",X"FF",X"77",X"27",X"72",X"27",X"70",X"70",X"27",X"72",X"27",X"77",X"FF",X"07",X"F0",
		X"0F",X"E0",X"FF",X"77",X"27",X"77",X"20",X"70",X"70",X"20",X"77",X"27",X"77",X"FF",X"E0",X"0F",
		X"00",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"E0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E7",X"E7",X"81",X"81",X"E7",X"E7",X"FF",
		X"01",X"03",X"01",X"01",X"07",X"03",X"01",X"03",X"1F",X"03",X"1F",X"0F",X"07",X"1F",X"03",X"0F",
		X"7F",X"0F",X"7F",X"3F",X"0F",X"7F",X"1F",X"3F",X"FF",X"3F",X"7F",X"FF",X"3F",X"FF",X"3F",X"7F",
		X"C4",X"CE",X"C4",X"CE",X"C0",X"C0",X"C0",X"C0",X"00",X"FF",X"FF",X"CE",X"C4",X"CE",X"C4",X"CE",
		X"CE",X"C4",X"CE",X"C4",X"CE",X"FF",X"FF",X"00",X"C0",X"C0",X"C0",X"C0",X"CE",X"C4",X"CE",X"C4",
		X"F0",X"07",X"FF",X"CE",X"C4",X"CE",X"C4",X"CE",X"0E",X"04",X"0E",X"04",X"0E",X"FF",X"07",X"F0",
		X"0F",X"E0",X"FF",X"CE",X"C4",X"CE",X"C4",X"CE",X"CE",X"C4",X"CE",X"C4",X"CE",X"FF",X"E0",X"0F",
		X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"E0",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"FF",X"E7",X"E7",X"FF",X"FF",X"E7",X"E7",X"FF",
		X"FF",X"FF",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"C3",X"C3",X"FF",X"FF",X"C3",X"C3",X"FF",X"00",X"00",X"00",X"00",X"FF",X"C3",X"C3",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"C3",X"FF",X"2F",X"03",X"3F",X"4F",X"FF",X"C3",X"C3",X"FF",
		X"FF",X"C3",X"C3",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"2F",X"03",X"3F",X"4F",X"00",X"00",X"00",X"00",
		X"FF",X"C3",X"C3",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"2F",X"03",X"3F",X"4F",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"C3",X"C3",X"FF",X"2F",X"03",X"3F",X"4F",X"00",X"00",X"00",X"00",X"2F",X"03",X"3F",X"4F",
		X"FF",X"FF",X"FF",X"FF",X"2F",X"03",X"3F",X"4F",X"2F",X"03",X"3F",X"4F",X"2F",X"03",X"3F",X"4F",
		X"9E",X"F2",X"F0",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"F0",X"F2",X"9E",
		X"9C",X"96",X"F2",X"F0",X"F0",X"F0",X"60",X"00",X"00",X"60",X"F0",X"F0",X"F0",X"F2",X"96",X"9C",
		X"F0",X"98",X"9C",X"F6",X"F2",X"F0",X"60",X"00",X"00",X"60",X"F0",X"F2",X"F6",X"9C",X"98",X"F0",
		X"F0",X"98",X"9C",X"F6",X"F2",X"62",X"00",X"00",X"00",X"62",X"F2",X"F6",X"9C",X"90",X"F0",X"F0",
		X"07",X"0C",X"38",X"60",X"C6",X"6C",X"38",X"00",X"00",X"38",X"6C",X"C6",X"60",X"38",X"0C",X"07",
		X"07",X"1C",X"70",X"C0",X"80",X"D8",X"70",X"00",X"00",X"70",X"D8",X"80",X"C0",X"70",X"1C",X"07",
		X"07",X"1C",X"70",X"C0",X"80",X"C0",X"60",X"00",X"00",X"60",X"C0",X"80",X"C0",X"70",X"1C",X"07",
		X"07",X"3C",X"60",X"C0",X"80",X"80",X"80",X"00",X"FF",X"80",X"80",X"80",X"C0",X"60",X"3C",X"0F",
		X"F8",X"FC",X"FC",X"FC",X"78",X"30",X"00",X"00",X"F8",X"7C",X"FE",X"FF",X"FF",X"FF",X"FE",X"F8",
		X"00",X"00",X"60",X"F8",X"FC",X"FC",X"F8",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7E",X"3C",
		X"78",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"1E",X"3F",X"7F",X"7F",X"3D",X"18",X"00",X"00",
		X"3F",X"7F",X"FF",X"FF",X"7F",X"3F",X"3F",X"1F",X"00",X"00",X"04",X"0E",X"1F",X"3F",X"3F",X"1F",
		X"00",X"80",X"C0",X"E0",X"E0",X"C0",X"C0",X"00",X"FF",X"7E",X"7C",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FE",X"00",X"03",X"07",X"0F",X"0F",X"0F",X"03",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"38",X"6C",X"7C",X"6C",X"38",X"00",X"38",X"6C",X"7C",X"6C",X"38",X"00",X"00",
		X"6C",X"7C",X"6C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",
		X"6C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"6C",X"7C",
		X"00",X"38",X"7C",X"E6",X"FE",X"E6",X"7C",X"38",X"7C",X"E6",X"FE",X"E6",X"7C",X"38",X"00",X"00",
		X"FE",X"E6",X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"E6",
		X"7C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"7C",X"E6",X"FE",X"E6",
		X"3C",X"7E",X"E7",X"FF",X"FF",X"E7",X"7E",X"3C",X"E7",X"FF",X"FF",X"E7",X"7E",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"7E",X"FF",X"E7",X"7E",X"3C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"3C",X"7E",X"E7",X"FF",X"7E",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"3C",X"7E",X"E7",X"FF",X"FF",X"E7",X"FF",X"CF",X"CE",X"FE",X"FC",X"70",X"00",X"00",
		X"00",X"00",X"00",X"70",X"FC",X"FE",X"CE",X"CF",X"07",X"07",X"03",X"03",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"FF",X"CF",X"CE",X"FE",X"FC",X"F8",X"F0",X"00",
		X"00",X"00",X"F0",X"F8",X"FC",X"FE",X"CE",X"CF",X"0E",X"0F",X"07",X"1F",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"03",X"1F",X"07",X"0F",X"7F",X"CE",X"CC",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"F8",X"CC",X"CE",X"1E",X"0F",X"27",X"3F",X"03",X"03",X"01",X"00",
		X"00",X"01",X"01",X"03",X"03",X"3F",X"27",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"27",X"33",X"1F",X"03",X"01",X"03",X"01",X"03",X"03",X"01",X"07",X"03",X"3F",X"67",X"4F",
		X"0C",X"67",X"73",X"1F",X"01",X"00",X"07",X"03",X"07",X"0F",X"01",X"03",X"00",X"1F",X"73",X"67",
		X"4C",X"F8",X"F8",X"F0",X"F8",X"F0",X"E0",X"C0",X"F8",X"F0",X"F8",X"F8",X"4C",X"4E",X"7E",X"4E",
		X"73",X"1F",X"71",X"01",X"07",X"03",X"1F",X"0F",X"01",X"03",X"71",X"1F",X"73",X"06",X"0C",X"06",
		X"F8",X"F0",X"F8",X"F8",X"F0",X"E0",X"80",X"00",X"F8",X"F8",X"4C",X"4E",X"7F",X"4E",X"4C",X"F8",
		X"00",X"00",X"80",X"E0",X"F0",X"F8",X"F8",X"F0",X"31",X"60",X"07",X"03",X"07",X"1F",X"7F",X"FE",
		X"31",X"1F",X"32",X"64",X"08",X"64",X"32",X"1F",X"00",X"FE",X"7F",X"1F",X"07",X"1F",X"01",X"63",
		X"F8",X"F0",X"F0",X"E0",X"80",X"00",X"00",X"00",X"4C",X"4E",X"7F",X"4E",X"4C",X"F8",X"F8",X"F0",
		X"C0",X"E0",X"F0",X"F0",X"F8",X"F0",X"F8",X"F8",X"07",X"03",X"0F",X"07",X"1F",X"7E",X"F0",X"00",
		X"73",X"06",X"0C",X"06",X"73",X"1F",X"71",X"00",X"1F",X"7F",X"07",X"0F",X"01",X"03",X"71",X"1F",
		X"FE",X"9C",X"98",X"F0",X"F8",X"FC",X"FC",X"7E",X"3E",X"7E",X"FC",X"FC",X"F8",X"F0",X"98",X"9C",
		X"30",X"18",X"0C",X"1F",X"F7",X"61",X"C0",X"00",X"00",X"00",X"C0",X"61",X"F7",X"1F",X"0C",X"18",
		X"98",X"F0",X"F8",X"FC",X"FC",X"7E",X"3E",X"3E",X"FC",X"FC",X"F8",X"F0",X"98",X"9C",X"FE",X"9C",
		X"0D",X"1F",X"FB",X"31",X"E0",X"00",X"00",X"00",X"E0",X"31",X"FB",X"1F",X"0D",X"19",X"31",X"19",
		X"F8",X"FC",X"FC",X"7E",X"3E",X"7F",X"1F",X"3F",X"F8",X"F0",X"98",X"9C",X"FE",X"9C",X"98",X"F0",
		X"3F",X"0F",X"1F",X"3F",X"3E",X"7E",X"FC",X"FC",X"3B",X"F1",X"20",X"E0",X"00",X"00",X"00",X"00",
		X"3B",X"1F",X"0D",X"19",X"39",X"19",X"0D",X"1F",X"00",X"00",X"00",X"00",X"00",X"E0",X"20",X"F1",
		X"FC",X"7E",X"3E",X"7F",X"1F",X"7F",X"1F",X"3F",X"98",X"9C",X"FE",X"9C",X"98",X"F0",X"F8",X"FC",
		X"3F",X"1F",X"7E",X"7E",X"FC",X"FC",X"F8",X"F0",X"0D",X"19",X"31",X"19",X"0D",X"EF",X"3B",X"E1",
		X"00",X"00",X"00",X"00",X"00",X"E1",X"3B",X"EF",X"7F",X"4E",X"CC",X"F8",X"F8",X"FC",X"FC",X"7C",
		X"FC",X"FC",X"FC",X"7C",X"F8",X"F8",X"CC",X"4E",X"0C",X"06",X"63",X"3F",X"61",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"61",X"3F",X"63",X"06",X"98",X"F0",X"F8",X"FC",X"FC",X"00",X"00",X"00",
		X"F8",X"FC",X"FC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"F8",
		X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",
		X"07",X"0F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"0F",
		X"0F",X"07",X"1F",X"7E",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"7E",X"0F",X"3F",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"3F",X"7E",X"F8",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F8",X"7E",X"0F",X"3F",X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"7F",
		X"1F",X"0F",X"1E",X"0E",X"1E",X"0C",X"1C",X"18",X"7E",X"3F",X"FF",X"1F",X"3F",X"0F",X"3F",X"0F",
		X"3F",X"0F",X"07",X"1F",X"0F",X"3F",X"1F",X"7E",X"00",X"18",X"1C",X"0C",X"1E",X"0E",X"1E",X"0F",
		X"1E",X"0E",X"3C",X"1C",X"18",X"30",X"00",X"00",X"70",X"38",X"3C",X"1C",X"3E",X"0E",X"3F",X"0F",
		X"0E",X"1E",X"1C",X"38",X"30",X"00",X"00",X"00",X"0F",X"3F",X"0F",X"3F",X"0F",X"1F",X"0E",X"1E",
		X"1F",X"0F",X"3F",X"0F",X"1F",X"0F",X"3F",X"0F",X"00",X"00",X"00",X"00",X"00",X"38",X"1C",X"0C",
		X"0E",X"1C",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"1C",X"0C",X"1E",X"0E",
		X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"FE",X"3E",X"7E",X"3C",X"7C",X"FC",X"78",X"F8",
		X"03",X"01",X"07",X"03",X"07",X"1E",X"00",X"00",X"F8",X"78",X"FC",X"7C",X"FC",X"3E",X"7E",X"3E",
		X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"00",X"00",X"00",X"1F",X"07",X"03",X"07",X"01",
		X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"C0",X"E0",X"F0",X"F8",X"F8",
		X"00",X"01",X"00",X"07",X"03",X"0F",X"1F",X"7C",X"00",X"7C",X"3F",X"0F",X"07",X"03",X"01",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		if(ce = '1') then data <= rom_data(to_integer(unsigned(addr))); end if;
	end if;
end process;
end architecture;
